module cex();

endmodule